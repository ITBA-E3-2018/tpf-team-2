module ToVGA (clk,hsync,vsync,r,g,b);
input wire clk;
output wire hsync,vsync,r,g,b;
parameter ADDRESS, FPORCH, BPORCH, HSYNC, VSYNC; //posicion de memoria donde arranca a estar guardada la pantalla que voy a mostrar.


endmodule