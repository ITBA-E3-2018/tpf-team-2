module mod1 (o, a, b);

input a,b;
output reg o;

and (o, a, b);

endmodule 